library verilog;
use verilog.vl_types.all;
entity \BUFFER\ is
    port(
        \OUT\           : out    vl_logic;
        \IN\            : in     vl_logic
    );
end \BUFFER\;
