module LCD_CTRL(clk, reset, IROM_Q, cmd, cmd_valid, IROM_EN, IROM_A, IRB_RW, IRB_D, IRB_A, busy, done);

input clk;
input reset;
input [7:0] IROM_Q;
input [2:0] cmd;
input cmd_valid;

output reg IROM_EN; // 0 for start to read, 1 for close IROM
output reg [5:0] IROM_A;
output reg IRB_RW;  // 0 for start to write, 1 for close IRB(?)
output reg [7:0] IRB_D;
output reg [5:0] IRB_A;
output reg busy;    // 1 for controller is executing current command, 0 for system to input the command, default is 1 when reseted
output reg done;    // 1 for controller finished writing to IRB

reg [2:0] curr_x, curr_y;
reg [3:0] curr_state, next_state;
reg [7:0] buffer [0:63];
//wire 		IROM_EN;
parameter Reset = 3'b000;
parameter Input = 3'b001;
//assign	IROM_EN = (curr_state==Input) ? 1'b0 : 1'b1;
always@(posedge clk) begin
    if(reset) begin
        
        busy <= 1;
        done <= 0;
        IRB_A <= 0;
        IRB_D <= 0;
        IRB_RW <= 1;
        curr_state <= Reset;
    end
    else begin
        curr_state <= next_state;
        case(curr_state) 
            Input: begin
               buffer[IROM_A] <= IROM_Q; 
            end
        endcase
    end
end

always@(*) begin
    //next_state = curr_state;
    case(curr_state) 
        Reset: begin
            next_state = Input;
            //IROM_EN <= 1;
            IROM_A = 63;
        end
        Input: begin
            IROM_A = (IROM_A == 63) ? 0 : IROM_A + 1;
            IROM_EN = (IROM_A == 63) ? 1 : 0;
            
            next_state = Input;

        end
    endcase
    

end

endmodule
