library verilog;
use verilog.vl_types.all;
entity CONV is
    generic(
        \WAIT\          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        LOAD            : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi1);
        NO_REUSE        : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi0);
        REUSE           : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi1, Hi1);
        CONVOLUTION_0   : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi0);
        RELU_0          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi0, Hi1);
        CONVOLUTION_1   : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi0);
        RELU_1          : vl_logic_vector(0 to 3) := (Hi0, Hi1, Hi1, Hi1);
        PRE_MAXPOOL     : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi0);
        MAXPOOL_0       : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi0, Hi1);
        MAXPOOL_1       : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi0);
        FLATTEN         : vl_logic_vector(0 to 3) := (Hi1, Hi0, Hi1, Hi1);
        ker0_0          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        ker0_1          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        ker0_2          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        ker0_3          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        ker0_4          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        ker0_5          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        ker0_6          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        ker0_7          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        ker0_8          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        ker1_0          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1);
        ker1_1          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0);
        ker1_2          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        ker1_3          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1);
        ker1_4          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        ker1_5          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1);
        ker1_6          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1);
        ker1_7          : vl_logic_vector(0 to 19) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        ker1_8          : vl_logic_vector(0 to 19) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        bias_0          : vl_logic_vector(0 to 39) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        bias_1          : vl_logic_vector(0 to 39) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0)
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        busy            : out    vl_logic;
        ready           : in     vl_logic;
        iaddr           : out    vl_logic_vector(11 downto 0);
        idata           : in     vl_logic_vector(19 downto 0);
        cwr             : out    vl_logic;
        caddr_wr        : out    vl_logic_vector(11 downto 0);
        cdata_wr        : out    vl_logic_vector(19 downto 0);
        crd             : out    vl_logic;
        caddr_rd        : out    vl_logic_vector(11 downto 0);
        cdata_rd        : in     vl_logic_vector(19 downto 0);
        csel            : out    vl_logic_vector(2 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of \WAIT\ : constant is 1;
    attribute mti_svvh_generic_type of LOAD : constant is 1;
    attribute mti_svvh_generic_type of NO_REUSE : constant is 1;
    attribute mti_svvh_generic_type of REUSE : constant is 1;
    attribute mti_svvh_generic_type of CONVOLUTION_0 : constant is 1;
    attribute mti_svvh_generic_type of RELU_0 : constant is 1;
    attribute mti_svvh_generic_type of CONVOLUTION_1 : constant is 1;
    attribute mti_svvh_generic_type of RELU_1 : constant is 1;
    attribute mti_svvh_generic_type of PRE_MAXPOOL : constant is 1;
    attribute mti_svvh_generic_type of MAXPOOL_0 : constant is 1;
    attribute mti_svvh_generic_type of MAXPOOL_1 : constant is 1;
    attribute mti_svvh_generic_type of FLATTEN : constant is 1;
    attribute mti_svvh_generic_type of ker0_0 : constant is 1;
    attribute mti_svvh_generic_type of ker0_1 : constant is 1;
    attribute mti_svvh_generic_type of ker0_2 : constant is 1;
    attribute mti_svvh_generic_type of ker0_3 : constant is 1;
    attribute mti_svvh_generic_type of ker0_4 : constant is 1;
    attribute mti_svvh_generic_type of ker0_5 : constant is 1;
    attribute mti_svvh_generic_type of ker0_6 : constant is 1;
    attribute mti_svvh_generic_type of ker0_7 : constant is 1;
    attribute mti_svvh_generic_type of ker0_8 : constant is 1;
    attribute mti_svvh_generic_type of ker1_0 : constant is 1;
    attribute mti_svvh_generic_type of ker1_1 : constant is 1;
    attribute mti_svvh_generic_type of ker1_2 : constant is 1;
    attribute mti_svvh_generic_type of ker1_3 : constant is 1;
    attribute mti_svvh_generic_type of ker1_4 : constant is 1;
    attribute mti_svvh_generic_type of ker1_5 : constant is 1;
    attribute mti_svvh_generic_type of ker1_6 : constant is 1;
    attribute mti_svvh_generic_type of ker1_7 : constant is 1;
    attribute mti_svvh_generic_type of ker1_8 : constant is 1;
    attribute mti_svvh_generic_type of bias_0 : constant is 1;
    attribute mti_svvh_generic_type of bias_1 : constant is 1;
end CONV;
