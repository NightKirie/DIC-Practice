library verilog;
use verilog.vl_types.all;
entity testfixture0 is
end testfixture0;
