module avg(din, reset, clk, ready, dout);
input reset, clk;
input [15:0] din;
output ready;
output [15:0] dout;

// ==========================================
//  Enter your design below
// ==========================================





endmodule
